`timescale 1ns/1ns

module And(
	input dato1,
	input dato2,
	output datoS
);

	assign datoS = dato1 & dato2;
endmodule
